Dot dot1 #(parameter x=13, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten1));
Dot dot2 #(parameter x=22, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten2));
Dot dot3 #(parameter x=31, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten3));
Dot dot4 #(parameter x=40, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten4));
Dot dot5 #(parameter x=49, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten5));
Dot dot6 #(parameter x=58, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten6));
Dot dot7 #(parameter x=67, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten7));
Dot dot8 #(parameter x=76, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten8));
Dot dot9 #(parameter x=85, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten9));
Dot dot10 #(parameter x=94, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten10));
Dot dot11 #(parameter x=103, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten11));
Dot dot12 #(parameter x=112, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten12));
Dot dot13 #(parameter x=140, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten13));
Dot dot14 #(parameter x=149, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten14));
Dot dot15 #(parameter x=158, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten15));
Dot dot16 #(parameter x=167, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten16));
Dot dot17 #(parameter x=176, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten17));
Dot dot18 #(parameter x=185, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten18));
Dot dot19 #(parameter x=194, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten19));
Dot dot20 #(parameter x=203, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten20));
Dot dot21 #(parameter x=212, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten21));
Dot dot22 #(parameter x=221, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten22));
Dot dot23 #(parameter x=230, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten23));
Dot dot24 #(parameter x=239, parameter y=10)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten24));
Dot dot25 #(parameter x=13, parameter y=19)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten25));
Dot dot26 #(parameter x=58, parameter y=19)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten26));
Dot dot27 #(parameter x=112, parameter y=19)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten27));
Dot dot28 #(parameter x=139, parameter y=19)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten28));
Dot dot29 #(parameter x=194, parameter y=19)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten29));
Dot dot30 #(parameter x=239, parameter y=19)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten30));
Dot dot31 #(parameter x=58, parameter y=27)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten31));
Dot dot32 #(parameter x=112, parameter y=27)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten32));
Dot dot33 #(parameter x=139, parameter y=27)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten33));
Dot dot34 #(parameter x=194, parameter y=27)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten34));
Dot dot35 #(parameter x=13, parameter y=35)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten35));
Dot dot36 #(parameter x=58, parameter y=35)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten36));
Dot dot37 #(parameter x=112, parameter y=35)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten37));
Dot dot38 #(parameter x=139, parameter y=35)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten38));
Dot dot39 #(parameter x=194, parameter y=35)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten39));
Dot dot40 #(parameter x=239, parameter y=35)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten40));
Dot dot41 #(parameter x=13, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten41));
Dot dot42 #(parameter x=22, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten42));
Dot dot43 #(parameter x=31, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten43));
Dot dot44 #(parameter x=40, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten44));
Dot dot45 #(parameter x=49, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten45));
Dot dot46 #(parameter x=58, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten46));
Dot dot47 #(parameter x=67, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten47));
Dot dot48 #(parameter x=76, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten48));
Dot dot49 #(parameter x=85, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten49));
Dot dot50 #(parameter x=95, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten50));
Dot dot51 #(parameter x=104, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten51));
Dot dot52 #(parameter x=113, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten52));
Dot dot53 #(parameter x=122, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten53));
Dot dot54 #(parameter x=131, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten54));
Dot dot55 #(parameter x=140, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten55));
Dot dot56 #(parameter x=149, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten56));
Dot dot57 #(parameter x=158, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten57));
Dot dot58 #(parameter x=167, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten58));
Dot dot59 #(parameter x=176, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten59));
Dot dot60 #(parameter x=185, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten60));
Dot dot61 #(parameter x=194, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten61));
Dot dot62 #(parameter x=203, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten62));
Dot dot63 #(parameter x=212, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten63));
Dot dot64 #(parameter x=221, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten64));
Dot dot65 #(parameter x=230, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten65));
Dot dot66 #(parameter x=240, parameter y=43)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten66));
Dot dot67 #(parameter x=13, parameter y=52)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten67));
Dot dot68 #(parameter x=58, parameter y=52)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten68));
Dot dot69 #(parameter x=85, parameter y=52)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten69));
Dot dot70 #(parameter x=167, parameter y=52)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten70));
Dot dot71 #(parameter x=194, parameter y=52)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten71));
Dot dot72 #(parameter x=239, parameter y=52)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten72));
Dot dot73 #(parameter x=13, parameter y=60)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten73));
Dot dot74 #(parameter x=58, parameter y=60)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten74));
Dot dot75 #(parameter x=85, parameter y=60)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten75));
Dot dot76 #(parameter x=167, parameter y=60)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten76));
Dot dot77 #(parameter x=194, parameter y=60)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten77));
Dot dot78 #(parameter x=239, parameter y=60)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten78));
Dot dot79 #(parameter x=13, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten79));
Dot dot80 #(parameter x=22, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten80));
Dot dot81 #(parameter x=31, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten81));
Dot dot82 #(parameter x=40, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten82));
Dot dot83 #(parameter x=49, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten83));
Dot dot84 #(parameter x=58, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten84));
Dot dot85 #(parameter x=85, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten85));
Dot dot86 #(parameter x=94, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten86));
Dot dot87 #(parameter x=103, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten87));
Dot dot88 #(parameter x=112, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten88));
Dot dot89 #(parameter x=139, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten89));
Dot dot90 #(parameter x=149, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten90));
Dot dot91 #(parameter x=158, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten91));
Dot dot92 #(parameter x=167, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten92));
Dot dot93 #(parameter x=194, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten93));
Dot dot94 #(parameter x=203, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten94));
Dot dot95 #(parameter x=212, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten95));
Dot dot96 #(parameter x=221, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten96));
Dot dot97 #(parameter x=230, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten97));
Dot dot98 #(parameter x=239, parameter y=68)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten98));
Dot dot99 #(parameter x=58, parameter y=76)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten99));
Dot dot100 #(parameter x=194, parameter y=76)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten100));
Dot dot101 #(parameter x=58, parameter y=85)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten101));
Dot dot102 #(parameter x=194, parameter y=85)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten102));
Dot dot103 #(parameter x=58, parameter y=93)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten103));
Dot dot104 #(parameter x=194, parameter y=93)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten104));
Dot dot105 #(parameter x=58, parameter y=101)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten105));
Dot dot106 #(parameter x=194, parameter y=101)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten106));
Dot dot107 #(parameter x=58, parameter y=110)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten107));
Dot dot108 #(parameter x=194, parameter y=110)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten108));
Dot dot109 #(parameter x=58, parameter y=118)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten109));
Dot dot110 #(parameter x=194, parameter y=118)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten110));
Dot dot111 #(parameter x=58, parameter y=126)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten111));
Dot dot112 #(parameter x=194, parameter y=126)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten112));
Dot dot113 #(parameter x=58, parameter y=134)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten113));
Dot dot114 #(parameter x=194, parameter y=134)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten114));
Dot dot115 #(parameter x=58, parameter y=143)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten115));
Dot dot116 #(parameter x=194, parameter y=143)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten116));
Dot dot117 #(parameter x=58, parameter y=151)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten117));
Dot dot118 #(parameter x=194, parameter y=151)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten118));
Dot dot119 #(parameter x=58, parameter y=159)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten119));
Dot dot120 #(parameter x=194, parameter y=159)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten120));
Dot dot121 #(parameter x=13, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten121));
Dot dot122 #(parameter x=22, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten122));
Dot dot123 #(parameter x=31, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten123));
Dot dot124 #(parameter x=40, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten124));
Dot dot125 #(parameter x=49, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten125));
Dot dot126 #(parameter x=58, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten126));
Dot dot127 #(parameter x=67, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten127));
Dot dot128 #(parameter x=76, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten128));
Dot dot129 #(parameter x=85, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten129));
Dot dot130 #(parameter x=94, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten130));
Dot dot131 #(parameter x=103, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten131));
Dot dot132 #(parameter x=112, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten132));
Dot dot133 #(parameter x=140, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten133));
Dot dot134 #(parameter x=149, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten134));
Dot dot135 #(parameter x=158, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten135));
Dot dot136 #(parameter x=167, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten136));
Dot dot137 #(parameter x=176, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten137));
Dot dot138 #(parameter x=185, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten138));
Dot dot139 #(parameter x=194, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten139));
Dot dot140 #(parameter x=203, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten140));
Dot dot141 #(parameter x=212, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten141));
Dot dot142 #(parameter x=221, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten142));
Dot dot143 #(parameter x=230, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten143));
Dot dot144 #(parameter x=239, parameter y=167)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten144));
Dot dot145 #(parameter x=13, parameter y=176)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten145));
Dot dot146 #(parameter x=58, parameter y=176)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten146));
Dot dot147 #(parameter x=112, parameter y=176)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten147));
Dot dot148 #(parameter x=139, parameter y=176)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten148));
Dot dot149 #(parameter x=194, parameter y=176)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten149));
Dot dot150 #(parameter x=239, parameter y=176)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten150));
Dot dot151 #(parameter x=13, parameter y=184)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten151));
Dot dot152 #(parameter x=58, parameter y=184)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten152));
Dot dot153 #(parameter x=112, parameter y=184)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten153));
Dot dot154 #(parameter x=139, parameter y=184)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten154));
Dot dot155 #(parameter x=194, parameter y=184)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten155));
Dot dot156 #(parameter x=239, parameter y=184)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten156));
Dot dot157 #(parameter x=22, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten157));
Dot dot158 #(parameter x=31, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten158));
Dot dot159 #(parameter x=58, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten159));
Dot dot160 #(parameter x=67, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten160));
Dot dot161 #(parameter x=76, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten161));
Dot dot162 #(parameter x=85, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten162));
Dot dot163 #(parameter x=94, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten163));
Dot dot164 #(parameter x=103, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten164));
Dot dot165 #(parameter x=112, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten165));
Dot dot166 #(parameter x=139, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten166));
Dot dot167 #(parameter x=148, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten167));
Dot dot168 #(parameter x=158, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten168));
Dot dot169 #(parameter x=167, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten169));
Dot dot170 #(parameter x=176, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten170));
Dot dot171 #(parameter x=185, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten171));
Dot dot172 #(parameter x=194, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten172));
Dot dot173 #(parameter x=221, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten173));
Dot dot174 #(parameter x=230, parameter y=192)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten174));
Dot dot175 #(parameter x=31, parameter y=200)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten175));
Dot dot176 #(parameter x=58, parameter y=200)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten176));
Dot dot177 #(parameter x=85, parameter y=200)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten177));
Dot dot178 #(parameter x=167, parameter y=200)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten178));
Dot dot179 #(parameter x=194, parameter y=200)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten179));
Dot dot180 #(parameter x=221, parameter y=200)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten180));
Dot dot181 #(parameter x=31, parameter y=209)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten181));
Dot dot182 #(parameter x=58, parameter y=209)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten182));
Dot dot183 #(parameter x=85, parameter y=209)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten183));
Dot dot184 #(parameter x=167, parameter y=209)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten184));
Dot dot185 #(parameter x=194, parameter y=209)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten185));
Dot dot186 #(parameter x=221, parameter y=209)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten186));
Dot dot187 #(parameter x=13, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten187));
Dot dot188 #(parameter x=22, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten188));
Dot dot189 #(parameter x=31, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten189));
Dot dot190 #(parameter x=40, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten190));
Dot dot191 #(parameter x=49, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten191));
Dot dot192 #(parameter x=58, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten192));
Dot dot193 #(parameter x=85, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten193));
Dot dot194 #(parameter x=94, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten194));
Dot dot195 #(parameter x=103, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten195));
Dot dot196 #(parameter x=112, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten196));
Dot dot197 #(parameter x=139, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten197));
Dot dot198 #(parameter x=148, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten198));
Dot dot199 #(parameter x=158, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten199));
Dot dot200 #(parameter x=167, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten200));
Dot dot201 #(parameter x=194, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten201));
Dot dot202 #(parameter x=203, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten202));
Dot dot203 #(parameter x=212, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten203));
Dot dot204 #(parameter x=221, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten204));
Dot dot205 #(parameter x=230, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten205));
Dot dot206 #(parameter x=239, parameter y=217)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten206));
Dot dot207 #(parameter x=13, parameter y=225)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten207));
Dot dot208 #(parameter x=112, parameter y=225)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten208));
Dot dot209 #(parameter x=139, parameter y=225)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten209));
Dot dot210 #(parameter x=239, parameter y=225)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten210));
Dot dot211 #(parameter x=13, parameter y=233)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten211));
Dot dot212 #(parameter x=112, parameter y=233)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten212));
Dot dot213 #(parameter x=140, parameter y=233)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten213));
Dot dot214 #(parameter x=239, parameter y=233)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten214));
Dot dot215 #(parameter x=13, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten215));
Dot dot216 #(parameter x=22, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten216));
Dot dot217 #(parameter x=31, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten217));
Dot dot218 #(parameter x=40, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten218));
Dot dot219 #(parameter x=49, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten219));
Dot dot220 #(parameter x=58, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten220));
Dot dot221 #(parameter x=67, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten221));
Dot dot222 #(parameter x=76, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten222));
Dot dot223 #(parameter x=85, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten223));
Dot dot224 #(parameter x=94, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten224));
Dot dot225 #(parameter x=103, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten225));
Dot dot226 #(parameter x=112, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten226));
Dot dot227 #(parameter x=121, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten227));
Dot dot228 #(parameter x=130, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten228));
Dot dot229 #(parameter x=139, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten229));
Dot dot230 #(parameter x=148, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten230));
Dot dot231 #(parameter x=158, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten231));
Dot dot232 #(parameter x=167, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten232));
Dot dot233 #(parameter x=176, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten233));
Dot dot234 #(parameter x=185, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten234));
Dot dot235 #(parameter x=194, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten235));
Dot dot236 #(parameter x=203, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten236));
Dot dot237 #(parameter x=212, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten237));
Dot dot238 #(parameter x=221, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten238));
Dot dot239 #(parameter x=230, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten239));
Dot dot240 #(parameter x=239, parameter y=242)(.Clk(CLK), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_X_Pos(pac_X_Pos), .pac_Y_Pos(pac_Y_Pos), .isEaten(isEaten240));

Dot #(13, 10) dot1 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten1));
Dot #(22, 10) dot2 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten2));
Dot #(31, 10) dot3 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten3));
Dot #(40, 10) dot4 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten4));
Dot #(49, 10) dot5 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten5));
Dot #(58, 10) dot6 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten6));
Dot #(67, 10) dot7 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten7));
Dot #(76, 10) dot8 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten8));
Dot #(85, 10) dot9 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten9));
Dot #(94, 10) dot10 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten10));
Dot #(103, 10) dot11 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten11));
Dot #(112, 10) dot12 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten12));
Dot #(140, 10) dot13 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten13));
Dot #(149, 10) dot14 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten14));
Dot #(158, 10) dot15 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten15));
Dot #(167, 10) dot16 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten16));
Dot #(176, 10) dot17 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten17));
Dot #(185, 10) dot18 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten18));
Dot #(194, 10) dot19 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten19));
Dot #(203, 10) dot20 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten20));
Dot #(212, 10) dot21 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten21));
Dot #(221, 10) dot22 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten22));
Dot #(230, 10) dot23 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten23));
Dot #(239, 10) dot24 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten24));
Dot #(13, 19) dot25 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten25));
Dot #(58, 19) dot26 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten26));
Dot #(112, 19) dot27 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten27));
Dot #(139, 19) dot28 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten28));
Dot #(194, 19) dot29 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten29));
Dot #(239, 19) dot30 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten30));
Dot #(58, 27) dot31 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten31));
Dot #(112, 27) dot32 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten32));
Dot #(139, 27) dot33 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten33));
Dot #(194, 27) dot34 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten34));
Dot #(13, 35) dot35 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten35));
Dot #(58, 35) dot36 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten36));
Dot #(112, 35) dot37 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten37));
Dot #(139, 35) dot38 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten38));
Dot #(194, 35) dot39 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten39));
Dot #(239, 35) dot40 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten40));
Dot #(13, 43) dot41 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten41));
Dot #(22, 43) dot42 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten42));
Dot #(31, 43) dot43 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten43));
Dot #(40, 43) dot44 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten44));
Dot #(49, 43) dot45 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten45));
Dot #(58, 43) dot46 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten46));
Dot #(67, 43) dot47 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten47));
Dot #(76, 43) dot48 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten48));
Dot #(85, 43) dot49 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten49));
Dot #(95, 43) dot50 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten50));
Dot #(104, 43) dot51 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten51));
Dot #(113, 43) dot52 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten52));
Dot #(122, 43) dot53 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten53));
Dot #(131, 43) dot54 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten54));
Dot #(140, 43) dot55 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten55));
Dot #(149, 43) dot56 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten56));
Dot #(158, 43) dot57 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten57));
Dot #(167, 43) dot58 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten58));
Dot #(176, 43) dot59 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten59));
Dot #(185, 43) dot60 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten60));
Dot #(194, 43) dot61 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten61));
Dot #(203, 43) dot62 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten62));
Dot #(212, 43) dot63 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten63));
Dot #(221, 43) dot64 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten64));
Dot #(230, 43) dot65 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten65));
Dot #(240, 43) dot66 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten66));
Dot #(13, 52) dot67 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten67));
Dot #(58, 52) dot68 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten68));
Dot #(85, 52) dot69 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten69));
Dot #(167, 52) dot70 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten70));
Dot #(194, 52) dot71 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten71));
Dot #(239, 52) dot72 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten72));
Dot #(13, 60) dot73 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten73));
Dot #(58, 60) dot74 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten74));
Dot #(85, 60) dot75 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten75));
Dot #(167, 60) dot76 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten76));
Dot #(194, 60) dot77 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten77));
Dot #(239, 60) dot78 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten78));
Dot #(13, 68) dot79 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten79));
Dot #(22, 68) dot80 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten80));
Dot #(31, 68) dot81 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten81));
Dot #(40, 68) dot82 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten82));
Dot #(49, 68) dot83 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten83));
Dot #(58, 68) dot84 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten84));
Dot #(85, 68) dot85 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten85));
Dot #(94, 68) dot86 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten86));
Dot #(103, 68) dot87 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten87));
Dot #(112, 68) dot88 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten88));
Dot #(139, 68) dot89 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten89));
Dot #(149, 68) dot90 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten90));
Dot #(158, 68) dot91 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten91));
Dot #(167, 68) dot92 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten92));
Dot #(194, 68) dot93 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten93));
Dot #(203, 68) dot94 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten94));
Dot #(212, 68) dot95 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten95));
Dot #(221, 68) dot96 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten96));
Dot #(230, 68) dot97 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten97));
Dot #(239, 68) dot98 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten98));
Dot #(58, 76) dot99 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten99));
Dot #(194, 76) dot100 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten100));
Dot #(58, 85) dot101 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten101));
Dot #(194, 85) dot102 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten102));
Dot #(58, 93) dot103 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten103));
Dot #(194, 93) dot104 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten104));
Dot #(58, 101) dot105 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten105));
Dot #(194, 101) dot106 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten106));
Dot #(58, 110) dot107 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten107));
Dot #(194, 110) dot108 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten108));
Dot #(58, 118) dot109 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten109));
Dot #(194, 118) dot110 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten110));
Dot #(58, 126) dot111 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten111));
Dot #(194, 126) dot112 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten112));
Dot #(58, 134) dot113 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten113));
Dot #(194, 134) dot114 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten114));
Dot #(58, 143) dot115 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten115));
Dot #(194, 143) dot116 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten116));
Dot #(58, 151) dot117 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten117));
Dot #(194, 151) dot118 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten118));
Dot #(58, 159) dot119 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten119));
Dot #(194, 159) dot120 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten120));
Dot #(13, 167) dot121 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten121));
Dot #(22, 167) dot122 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten122));
Dot #(31, 167) dot123 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten123));
Dot #(40, 167) dot124 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten124));
Dot #(49, 167) dot125 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten125));
Dot #(58, 167) dot126 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten126));
Dot #(67, 167) dot127 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten127));
Dot #(76, 167) dot128 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten128));
Dot #(85, 167) dot129 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten129));
Dot #(94, 167) dot130 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten130));
Dot #(103, 167) dot131 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten131));
Dot #(112, 167) dot132 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten132));
Dot #(140, 167) dot133 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten133));
Dot #(149, 167) dot134 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten134));
Dot #(158, 167) dot135 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten135));
Dot #(167, 167) dot136 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten136));
Dot #(176, 167) dot137 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten137));
Dot #(185, 167) dot138 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten138));
Dot #(194, 167) dot139 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten139));
Dot #(203, 167) dot140 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten140));
Dot #(212, 167) dot141 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten141));
Dot #(221, 167) dot142 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten142));
Dot #(230, 167) dot143 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten143));
Dot #(239, 167) dot144 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten144));
Dot #(13, 176) dot145 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten145));
Dot #(58, 176) dot146 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten146));
Dot #(112, 176) dot147 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten147));
Dot #(139, 176) dot148 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten148));
Dot #(194, 176) dot149 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten149));
Dot #(239, 176) dot150 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten150));
Dot #(13, 184) dot151 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten151));
Dot #(58, 184) dot152 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten152));
Dot #(112, 184) dot153 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten153));
Dot #(139, 184) dot154 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten154));
Dot #(194, 184) dot155 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten155));
Dot #(239, 184) dot156 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten156));
Dot #(22, 192) dot157 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten157));
Dot #(31, 192) dot158 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten158));
Dot #(58, 192) dot159 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten159));
Dot #(67, 192) dot160 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten160));
Dot #(76, 192) dot161 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten161));
Dot #(85, 192) dot162 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten162));
Dot #(94, 192) dot163 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten163));
Dot #(103, 192) dot164 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten164));
Dot #(112, 192) dot165 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten165));
Dot #(139, 192) dot166 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten166));
Dot #(148, 192) dot167 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten167));
Dot #(158, 192) dot168 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten168));
Dot #(167, 192) dot169 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten169));
Dot #(176, 192) dot170 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten170));
Dot #(185, 192) dot171 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten171));
Dot #(194, 192) dot172 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten172));
Dot #(221, 192) dot173 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten173));
Dot #(230, 192) dot174 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten174));
Dot #(31, 200) dot175 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten175));
Dot #(58, 200) dot176 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten176));
Dot #(85, 200) dot177 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten177));
Dot #(167, 200) dot178 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten178));
Dot #(194, 200) dot179 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten179));
Dot #(221, 200) dot180 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten180));
Dot #(31, 209) dot181 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten181));
Dot #(58, 209) dot182 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten182));
Dot #(85, 209) dot183 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten183));
Dot #(167, 209) dot184 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten184));
Dot #(194, 209) dot185 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten185));
Dot #(221, 209) dot186 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten186));
Dot #(13, 217) dot187 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten187));
Dot #(22, 217) dot188 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten188));
Dot #(31, 217) dot189 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten189));
Dot #(40, 217) dot190 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten190));
Dot #(49, 217) dot191 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten191));
Dot #(58, 217) dot192 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten192));
Dot #(85, 217) dot193 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten193));
Dot #(94, 217) dot194 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten194));
Dot #(103, 217) dot195 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten195));
Dot #(112, 217) dot196 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten196));
Dot #(139, 217) dot197 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten197));
Dot #(148, 217) dot198 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten198));
Dot #(158, 217) dot199 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten199));
Dot #(167, 217) dot200 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten200));
Dot #(194, 217) dot201 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten201));
Dot #(203, 217) dot202 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten202));
Dot #(212, 217) dot203 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten203));
Dot #(221, 217) dot204 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten204));
Dot #(230, 217) dot205 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten205));
Dot #(239, 217) dot206 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten206));
Dot #(13, 225) dot207 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten207));
Dot #(112, 225) dot208 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten208));
Dot #(139, 225) dot209 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten209));
Dot #(239, 225) dot210 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten210));
Dot #(13, 233) dot211 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten211));
Dot #(112, 233) dot212 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten212));
Dot #(140, 233) dot213 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten213));
Dot #(239, 233) dot214 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten214));
Dot #(13, 242) dot215 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten215));
Dot #(22, 242) dot216 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten216));
Dot #(31, 242) dot217 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten217));
Dot #(40, 242) dot218 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten218));
Dot #(49, 242) dot219 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten219));
Dot #(58, 242) dot220 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten220));
Dot #(67, 242) dot221 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten221));
Dot #(76, 242) dot222 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten222));
Dot #(85, 242) dot223 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten223));
Dot #(94, 242) dot224 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten224));
Dot #(103, 242) dot225 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten225));
Dot #(112, 242) dot226 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten226));
Dot #(121, 242) dot227 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten227));
Dot #(130, 242) dot228 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten228));
Dot #(139, 242) dot229 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten229));
Dot #(148, 242) dot230 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten230));
Dot #(158, 242) dot231 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten231));
Dot #(167, 242) dot232 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten232));
Dot #(176, 242) dot233 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten233));
Dot #(185, 242) dot234 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten234));
Dot #(194, 242) dot235 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten235));
Dot #(203, 242) dot236 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten236));
Dot #(212, 242) dot237 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten237));
Dot #(221, 242) dot238 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten238));
Dot #(230, 242) dot239 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten239));
Dot #(239, 242) dot240 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten240));

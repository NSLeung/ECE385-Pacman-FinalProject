//-------------------------------------------------------------------------
//      lab8.sv                                                          --
//      Christine Chen                                                   --
//      Fall 2014                                                        --
//                                                                       --
//      Modified by Po-Han Huang                                         --
//      10/06/2017                                                       --
//                                                                       --
//      Fall 2017 Distribution                                           --
//                                                                       --
//      For use with ECE 385 Lab 8                                       --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------


module final_top( input               CLOCK_50,
             input        [3:0]  KEY,          //bit 0 is set up as Reset
             output logic [6:0]  HEX0, HEX1,HEX2,HEX3,HEX4,HEX5,HEX6,HEX7,
             // VGA Interface
             output logic [7:0]  VGA_R,        //VGA Red
                                 VGA_G,        //VGA Green
                                 VGA_B,        //VGA Blue
             output logic        VGA_CLK,      //VGA Clock
                                 VGA_SYNC_N,   //VGA Sync signal
                                 VGA_BLANK_N,  //VGA Blank signal
                                 VGA_VS,       //VGA virtical sync signal
                                 VGA_HS,       //VGA horizontal sync signal
             // CY7C67200 Interface
             inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
             output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
             output logic        OTG_CS_N,     //CY7C67200 Chip Select
                                 OTG_RD_N,     //CY7C67200 Write
                                 OTG_WR_N,     //CY7C67200 Read
                                 OTG_RST_N,    //CY7C67200 Reset
             input               OTG_INT,      //CY7C67200 Interrupt
             // SDRAM Interface for Nios II Software
             output logic [12:0] DRAM_ADDR,    //SDRAM Address 13 Bits
             inout  wire  [31:0] DRAM_DQ,      //SDRAM Data 32 Bits
             output logic [1:0]  DRAM_BA,      //SDRAM Bank Address 2 Bits
             output logic [3:0]  DRAM_DQM,     //SDRAM Data Mast 4 Bits
             output logic        DRAM_RAS_N,   //SDRAM Row Address Strobe
                                 DRAM_CAS_N,   //SDRAM Column Address Strobe
                                 DRAM_CKE,     //SDRAM Clock Enable
                                 DRAM_WE_N,    //SDRAM Write Enable
                                 DRAM_CS_N,    //SDRAM Chip Select
                                 DRAM_CLK      //SDRAM Clock



                                 // SRAM controls (may be missing a clk signal??)
//                      				output logic [19:0] SRAM_ADDR,	// SRAM Address 20 Bits
//                      				inout wire [15:0] SRAM_DQ,			// SRAM Data 16 Bits
//                      				output logic 	SRAM_CE_N,			// SRAM Chip Enable
//                      									SRAM_LB_N,			// SRAM Lower Byte Enable (?)
//                      									SRAM_OE_N,			// SRAM Output Enable(?)
//                      									SRAM_UB_N,			// SRAM Upper Byte Enable (?)
//                      									SRAM_WE_N			// SRAM Write Enable (?)
                    );

    logic Reset_h, Clk, Reset_ball_h;
    logic [7:0] keycode;

    //logic for sram ctrl module
    logic ready, enable;
    // logic [15:0] SRAM_DATA, toSRAM_ctrl_data;
    logic [9:0]  DrawX, DrawY;
	  logic [19:0] frontbuff_addr, backbuff_addr;
	  // this was not initialised last night
	  logic SRAM_WE_CTRL;
//    logic [7:0] pac_X_Pos, pac_Y_Pos;

//    assign enable = ~(VGA_BLANK_N | ~FD_write_request_n);  //set enable 0 when the VGA is trying to read, and the frame_drawer wants to write.
//    assign SRAM_WE_CTRL = VGA_BLANK_N | FD_write_request_n; //always read (1) when not blanking (1) and if not writing (1)




    assign Clk = CLOCK_50;

    //clk counter for slowing down clk
    // logic [31:0] clk_counter = 32'd0;
    // logic clear;
    always_ff @ (posedge Clk) begin
        Reset_h <= ~(KEY[0]);        // The push buttons are active low
		  Reset_pac_h <= ~(KEY[2]);
      score_in <= score_out;
      // clear <=0;
      // if(clk_counter == 32'h005F5E100 )
      // begin
      //   clear <= 1'd1;
      //   clk_counter <= 0;
      // end
      // else clk_counter <= clk_counter + 32'd1;
    end

    //HPI interface logic variables
    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w, hpi_cs, hpi_reset;

    //address calculations done inside draw_controller
    logic [19:0] pixel_address;
	   logic [19:0] address;

     //logic variables for draw_control and color_mapper
     logic [3:0] color_index;
		logic [3:0] memtest;

    //logic variables for pac_controller
    logic isPac;
    logic [7:0] pac_mem_start_X, pac_mem_start_Y;

    //logic variables for AI_controller
    logic isAI;
    logic [7:0] AI_mem_start_X, AI_mem_start_Y;
    //ram.sv
    logic [3:0] mem_bg [0:65535];

    //scoreboard
    logic[7:0] score_out;
    logic[7:0] score_in = 8'b0;

    // always_ff @ (posedge VGA_VS)
    // begin
    //
    // end
    // Dot dot(score_in(score_in), score_out(score))
    //always comb block
    always_comb
    begin
      //initialize toSRAM_ctrl_data
      // toSRAM_ctrl_data = frontbuff_data;
      //address index into SRAM (pay attention width)
      //CHANGE HERE
//     pixel_address = DrawY_in * 19'd640 + DrawX_in;
		// pixel_address = DrawY_in * 19'd226 + DrawX_in; // Width of image is 226
    //  if (SRAM_WE_CTRL == 1'b1)
    //    address = pixel_address;
    //  else
			// address = 19'd0; // commented the next line because frontbuff is populated in the framebuffer module and this is the game logic which is not required for just the background.
      // address = frontbuff_addr;
    end

    // Interface between NIOS II and EZ-OTG chip
   hpi_io_intf hpi_io_inst(
                           .Clk(Clk),
                           .Reset(Reset_h),
                           // signals connected to NIOS II
                           .from_sw_address(hpi_addr),
                           .from_sw_data_in(hpi_data_in),
                           .from_sw_data_out(hpi_data_out),
                           .from_sw_r(hpi_r),
                           .from_sw_w(hpi_w),
                           .from_sw_cs(hpi_cs),
                           .from_sw_reset(hpi_reset),
                           // signals connected to EZ-OTG chip
                           .OTG_DATA(OTG_DATA),
                           .OTG_ADDR(OTG_ADDR),
                           .OTG_RD_N(OTG_RD_N),
                           .OTG_WR_N(OTG_WR_N),
                           .OTG_CS_N(OTG_CS_N),
                           .OTG_RST_N(OTG_RST_N)
   );
//
//     // You need to make sure that the port names here match the ports in Qsys-generated codes.
    pacman_finalproject_wkeycode_soc nios_system(
                            .clk_clk(Clk),
                            .reset_reset_n(1'b1),    // Never reset NIOS
                            .sdram_wire_addr(DRAM_ADDR),
                            .sdram_wire_ba(DRAM_BA),
                            .sdram_wire_cas_n(DRAM_CAS_N),
                            .sdram_wire_cke(DRAM_CKE),
                            .sdram_wire_cs_n(DRAM_CS_N),
                            .sdram_wire_dq(DRAM_DQ),
                            .sdram_wire_dqm(DRAM_DQM),
                            .sdram_wire_ras_n(DRAM_RAS_N),
                            .sdram_wire_we_n(DRAM_WE_N),
                            .sdram_clk_clk(DRAM_CLK),
                            .keycode_export(keycode),
                            .otg_hpi_address_export(hpi_addr),
                            .otg_hpi_data_in_port(hpi_data_in),
                            .otg_hpi_data_out_port(hpi_data_out),
                            .otg_hpi_cs_export(hpi_cs),
                            .otg_hpi_r_export(hpi_r),
                            .otg_hpi_w_export(hpi_w),
                            .otg_hpi_reset_export(hpi_reset)
   );

    // Use PLL to generate the 25MHZ VGA_CLK.
    // You will have to generate it on your own in simulation.
    vga_clk vga_clk_instance(.inclk0(Clk), .c0(VGA_CLK));
    // vga_clk vga_clk_instance(.inclk0(clear), .c0(VGA_CLK));


    // VGA Controller module
    // VGA_controller vga_controller_instance(.*, .Reset(Reset_h));
    VGA_controller vga_controller_instance(
                            .Reset(Reset_h),
                            .VGA_HS(VGA_HS),
                            .VGA_VS(VGA_VS),
                            .VGA_CLK(VGA_CLK),
                            .VGA_BLANK_N(VGA_BLANK_N),
                            .VGA_SYNC_N(VGA_SYNC_N),

                            //outputs from vga controller
                            .DrawX(DrawX),
														 .DrawY(DrawY)
    );

    // Which signal should be frame_clk?
    // ball ball_instance(.Clk(Clk), .Reset(Reset_ball_h), .frame_clk(VGA_VS), .DrawX(DrawX), .DrawY(DrawY), .keycode(keycode), .is_ball(is_ball));



    //color mapper module
    // color_mapper color_instance(.*);
    color_mapper color_instance(
                      //input
                        .color_index(color_index),


                        //output
                        .VGA_R(VGA_R),
                        .VGA_G(VGA_G),
                        .VGA_B(VGA_B)
    );

    //instantiate sram_ctrl
    // sram_ctrl sram_ctrl_module(
    //                   .clk(Clk),
    //                   .reset_n(~Reset_h),
    //                   .start_n(enable),
    //                   .addr_in(address),
    //                   .data_write(toSRAM_ctrl_data),
    //                   .rw(SRAM_WE_CTRL),  // 1  means read, 0 means write
    //                   //outputs
    //                   .ready(ready),
    //                   .data_read(SRAM_DATA),
    //                   .sram_addr(SRAM_ADDR),
    //                   .we_n(SRAM_WE_N),
    //                   .oe_n(SRAM_OE_N),
    //                   .ce_a_n(SRAM_CE_N),
    //                   .ub_a_n(SRAM_UB_N),
    //                   .lb_a_n(SRAM_LB_N),
    //                   .data_io(SRAM_DQ)
    // );

	 // Commented out frame_drawer for now because it determines the logic and position for the smaller sprites (Trying to get just the background now)
	 /*
    frame_drawer frame_drawer_instance(.CLK(Clk),
													.RESET(Reset_h),
													.ENABLE(VGA_BLANK_N),
													.DRAW_READY(ready),
                          //output
													.WRITEADDR(frontbuff_addr),


                          //COMING FROM SOFTWARE - NOT IMPLEMENTING YET
													// .PLAYER_X(player_coords[15:8]),
													// .PLAYER_Y(player_coords[7:0]),
													// .PLAYER_DIR(player_info[1:0]),
													.UI_ENABLE(1'b1),
													.DATA(fd_data),
													.DRAW_COMMAND(~KEY[3] | player_info[2]),
													.MAP_ID(player_info[6:4]),
													.FD_WE_N(FD_write_request_n),
													.ocm_data_out(temp_data)
    );

*/
    draw_control draw_control_instance(
                  .CLK(Clk),
                  // .CLK(clear),
                  .RESET(Reset_h),
                  // .ENABLE(VGA_BLANK_N),  //blanking enable for drawing
                  // .DRAW_READY(sram_done),

                  //input
                  .isPac(isPac),
                  .isAI(isAI),
						.isEaten(isEaten),
      				.DrawX(DrawX),
      				.DrawY(DrawY),
              .score_in(score_in),
              .score_out(score_out),
                  .pac_mem_start_X(pac_mem_start_X),
                  .pac_mem_start_Y(pac_mem_start_Y),
                  .AI_mem_start_X(AI_mem_start_X),
                  .AI_mem_start_Y(AI_mem_start_Y),
                  //outputs from draw_control
                   // .WRITEADDR(frontbuff_addr),
                   // .DATA(frontbuff_data),
                  // .FD_WE_N(FD_write_request_n),
                   .mem_address_out(address)
    );

    //Maze background here
    frameRAM frameRAM_instance(
    										// .write_address(16'b0), //don't care
    										.read_address(address),
    										.we(1'b0), //we always low

                        //input
                        .isPac(isPac),
                        .isAI(isAI),
    										.Clk(Clk),
    										.data_out(color_index)
                        ,.memdata(memtest),
                        .mem_bg(mem_bg)
    );

//		logic frame_clk_rising_edge;
    //instantiate pac module - determines whether pacman should be drawn or not
    pac_controller pacman(
          .Clk(CLK),
          // .Clk(clear),
          // .Reset(Reset_h),
          .Reset(Reset_pac_h),
          .frame_clk(VGA_VS),
          //raw_input
          .DrawX(DrawX),
          .DrawY(DrawY),
          .keycode(keycode),
//          .mem1(mem_bg),
          //hardcode keycode to enter default state
          // .keycode(8'h1F),
          .pac_mem_start_X(pac_mem_start_X),
          .pac_mem_start_Y(pac_mem_start_Y),
//          .pac_X_Pos(pac_X_Pos),
//          .pac_Y_Pos(pac_Y_Pos),
          //output
          .isPac(isPac)
    );

    AI_controller ai(
          .Clk(CLK),
          // .Clk(clear),
          // .Reset(Reset_h),
          .Reset(Reset_pac_h),
          .frame_clk(VGA_VS),
          //raw_input
          .DrawX(DrawX),
          .DrawY(DrawY),
          .AI_mem_start_X(AI_mem_start_X),
          .AI_mem_start_Y(AI_mem_start_Y),
          //output
          .isAI(isAI)
    );




    // Display keycode on hex display
    HexDriver hex_inst_0 ({2'b0, color_index[1:0]}, HEX0);
    HexDriver hex_inst_1 (keycode[3:0], HEX1);
    // HexDriver hex_inst_1 (DrawX[3:0], HEX1);
	 HexDriver hex_inst_2 (keycode[7:4], HEX2);
	 HexDriver hex_inst_3 (memtest, HEX3);
//	 HexDriver hex_inst_7 (frame_clk_rising_edge, HEX7);

   HexDriver hex_inst_4 (score_out[3:0], HEX4);
   HexDriver hex_inst_5 (score_out[7:4], HEX5);
   // HexDriver hex_inst_6 (score_out[11:8], HEX6);
   // HexDriver hex_inst_7 (clk_counter[14:11], HEX7);

assign isEaten = isEaten1 || isEaten2 || isEaten3 || isEaten4 || isEaten5 || isEaten6 || isEaten7 || isEaten8 || isEaten9 || isEaten10 || isEaten11 || isEaten12 || isEaten13 || isEaten14 || isEaten15 || isEaten16 || isEaten17 || isEaten18 || isEaten19 || isEaten20 || isEaten21 || isEaten22 || isEaten23 || isEaten24 || isEaten25 || isEaten26 || isEaten27 || isEaten28 || isEaten29 || isEaten30 || isEaten31 || isEaten32 || isEaten33 || isEaten34 || isEaten35 || isEaten36 || isEaten37 || isEaten38 || isEaten39 || isEaten40 || isEaten41 || isEaten42 || isEaten43 || isEaten44 || isEaten45 || isEaten46 || isEaten47 || isEaten48 || isEaten49 || isEaten50 || isEaten51 || isEaten52 || isEaten53 || isEaten54 || isEaten55 || isEaten56 || isEaten57 || isEaten58 || isEaten59 || isEaten60 || isEaten61 || isEaten62 || isEaten63 || isEaten64 || isEaten65 || isEaten66 || isEaten67 || isEaten68 || isEaten69 || isEaten70 || isEaten71 || isEaten72 || isEaten73 || isEaten74 || isEaten75 || isEaten76 || isEaten77 || isEaten78 || isEaten79 || isEaten80 || isEaten81 || isEaten82 || isEaten83 || isEaten84 || isEaten85 || isEaten86 || isEaten87 || isEaten88 || isEaten89 || isEaten90 || isEaten91 || isEaten92 || isEaten93 || isEaten94 || isEaten95 || isEaten96 || isEaten97 || isEaten98 || isEaten99 || isEaten100 || isEaten101 || isEaten102 || isEaten103 || isEaten104 || isEaten105 || isEaten106 || isEaten107 || isEaten108 || isEaten109 || isEaten110 || isEaten111 || isEaten112 || isEaten113 || isEaten114 || isEaten115 || isEaten116 || isEaten117 || isEaten118 || isEaten119 || isEaten120 || isEaten121 || isEaten122 || isEaten123 || isEaten124 || isEaten125 || isEaten126 || isEaten127 || isEaten128 || isEaten129 || isEaten130 || isEaten131 || isEaten132 || isEaten133 || isEaten134 || isEaten135 || isEaten136 || isEaten137 || isEaten138 || isEaten139 || isEaten140 || isEaten141 || isEaten142 || isEaten143 || isEaten144 || isEaten145 || isEaten146 || isEaten147 || isEaten148 || isEaten149 || isEaten150 || isEaten151 || isEaten152 || isEaten153 || isEaten154 || isEaten155 || isEaten156 || isEaten157 || isEaten158 || isEaten159 || isEaten160 || isEaten161 || isEaten162 || isEaten163 || isEaten164 || isEaten165 || isEaten166 || isEaten167 || isEaten168 || isEaten169 || isEaten170 || isEaten171 || isEaten172 || isEaten173 || isEaten174 || isEaten175 || isEaten176 || isEaten177 || isEaten178 || isEaten179 || isEaten180 || isEaten181 || isEaten182 || isEaten183 || isEaten184 || isEaten185 || isEaten186 || isEaten187 || isEaten188 || isEaten189 || isEaten190 || isEaten191 || isEaten192 || isEaten193 || isEaten194 || isEaten195 || isEaten196 || isEaten197 || isEaten198 || isEaten199 || isEaten200 || isEaten201 || isEaten202 || isEaten203 || isEaten204 || isEaten205 || isEaten206 || isEaten207 || isEaten208 || isEaten209 || isEaten210 || isEaten211 || isEaten212 || isEaten213 || isEaten214 || isEaten215 || isEaten216 || isEaten217 || isEaten218 || isEaten219 || isEaten220 || isEaten221 || isEaten222 || isEaten223 || isEaten224 || isEaten225 || isEaten226 || isEaten227 || isEaten228 || isEaten229 || isEaten230 || isEaten231 || isEaten232 || isEaten233 || isEaten234 || isEaten235 || isEaten236 || isEaten237 || isEaten238 || isEaten239 || isEaten240;


logic isEaten;

logic isEaten1;

logic isEaten2;

logic isEaten3;

logic isEaten4;

logic isEaten5;

logic isEaten6;

logic isEaten7;

logic isEaten8;

logic isEaten9;

logic isEaten10;

logic isEaten11;

logic isEaten12;

logic isEaten13;

logic isEaten14;

logic isEaten15;

logic isEaten16;

logic isEaten17;

logic isEaten18;

logic isEaten19;

logic isEaten20;

logic isEaten21;

logic isEaten22;

logic isEaten23;

logic isEaten24;

logic isEaten25;

logic isEaten26;

logic isEaten27;

logic isEaten28;

logic isEaten29;

logic isEaten30;

logic isEaten31;

logic isEaten32;

logic isEaten33;

logic isEaten34;

logic isEaten35;

logic isEaten36;

logic isEaten37;

logic isEaten38;

logic isEaten39;

logic isEaten40;

logic isEaten41;

logic isEaten42;

logic isEaten43;

logic isEaten44;

logic isEaten45;

logic isEaten46;

logic isEaten47;

logic isEaten48;

logic isEaten49;

logic isEaten50;

logic isEaten51;

logic isEaten52;

logic isEaten53;

logic isEaten54;

logic isEaten55;

logic isEaten56;

logic isEaten57;

logic isEaten58;

logic isEaten59;

logic isEaten60;

logic isEaten61;

logic isEaten62;

logic isEaten63;

logic isEaten64;

logic isEaten65;

logic isEaten66;

logic isEaten67;

logic isEaten68;

logic isEaten69;

logic isEaten70;

logic isEaten71;

logic isEaten72;

logic isEaten73;

logic isEaten74;

logic isEaten75;

logic isEaten76;

logic isEaten77;

logic isEaten78;

logic isEaten79;

logic isEaten80;

logic isEaten81;

logic isEaten82;

logic isEaten83;

logic isEaten84;

logic isEaten85;

logic isEaten86;

logic isEaten87;

logic isEaten88;

logic isEaten89;

logic isEaten90;

logic isEaten91;

logic isEaten92;

logic isEaten93;

logic isEaten94;

logic isEaten95;

logic isEaten96;

logic isEaten97;

logic isEaten98;

logic isEaten99;

logic isEaten100;

logic isEaten101;

logic isEaten102;

logic isEaten103;

logic isEaten104;

logic isEaten105;

logic isEaten106;

logic isEaten107;

logic isEaten108;

logic isEaten109;

logic isEaten110;

logic isEaten111;

logic isEaten112;

logic isEaten113;

logic isEaten114;

logic isEaten115;

logic isEaten116;

logic isEaten117;

logic isEaten118;

logic isEaten119;

logic isEaten120;

logic isEaten121;

logic isEaten122;

logic isEaten123;

logic isEaten124;

logic isEaten125;

logic isEaten126;

logic isEaten127;

logic isEaten128;

logic isEaten129;

logic isEaten130;

logic isEaten131;

logic isEaten132;

logic isEaten133;

logic isEaten134;

logic isEaten135;

logic isEaten136;

logic isEaten137;

logic isEaten138;

logic isEaten139;

logic isEaten140;

logic isEaten141;

logic isEaten142;

logic isEaten143;

logic isEaten144;

logic isEaten145;

logic isEaten146;

logic isEaten147;

logic isEaten148;

logic isEaten149;

logic isEaten150;

logic isEaten151;

logic isEaten152;

logic isEaten153;

logic isEaten154;

logic isEaten155;

logic isEaten156;

logic isEaten157;

logic isEaten158;

logic isEaten159;

logic isEaten160;

logic isEaten161;

logic isEaten162;

logic isEaten163;

logic isEaten164;

logic isEaten165;

logic isEaten166;

logic isEaten167;

logic isEaten168;

logic isEaten169;

logic isEaten170;

logic isEaten171;

logic isEaten172;

logic isEaten173;

logic isEaten174;

logic isEaten175;

logic isEaten176;

logic isEaten177;

logic isEaten178;

logic isEaten179;

logic isEaten180;

logic isEaten181;

logic isEaten182;

logic isEaten183;

logic isEaten184;

logic isEaten185;

logic isEaten186;

logic isEaten187;

logic isEaten188;

logic isEaten189;

logic isEaten190;

logic isEaten191;

logic isEaten192;

logic isEaten193;

logic isEaten194;

logic isEaten195;

logic isEaten196;

logic isEaten197;

logic isEaten198;

logic isEaten199;

logic isEaten200;

logic isEaten201;

logic isEaten202;

logic isEaten203;

logic isEaten204;

logic isEaten205;

logic isEaten206;

logic isEaten207;

logic isEaten208;

logic isEaten209;

logic isEaten210;

logic isEaten211;

logic isEaten212;

logic isEaten213;

logic isEaten214;

logic isEaten215;

logic isEaten216;

logic isEaten217;

logic isEaten218;

logic isEaten219;

logic isEaten220;

logic isEaten221;

logic isEaten222;

logic isEaten223;

logic isEaten224;

logic isEaten225;

logic isEaten226;

logic isEaten227;

logic isEaten228;

logic isEaten229;

logic isEaten230;

logic isEaten231;

logic isEaten232;

logic isEaten233;

logic isEaten234;

logic isEaten235;

logic isEaten236;

logic isEaten237;

logic isEaten238;

logic isEaten239;

logic isEaten240;

Dot #(13, 10) dot1 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten1));
Dot #(22, 10) dot2 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten2));
Dot #(31, 10) dot3 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten3));
Dot #(40, 10) dot4 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten4));
Dot #(49, 10) dot5 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten5));
Dot #(58, 10) dot6 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten6));
Dot #(67, 10) dot7 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten7));
Dot #(76, 10) dot8 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten8));
Dot #(85, 10) dot9 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten9));
Dot #(94, 10) dot10 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten10));
Dot #(103, 10) dot11 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten11));
Dot #(112, 10) dot12 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten12));
Dot #(140, 10) dot13 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten13));
Dot #(149, 10) dot14 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten14));
Dot #(158, 10) dot15 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten15));
Dot #(167, 10) dot16 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten16));
Dot #(176, 10) dot17 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten17));
Dot #(185, 10) dot18 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten18));
Dot #(194, 10) dot19 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten19));
Dot #(203, 10) dot20 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten20));
Dot #(212, 10) dot21 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten21));
Dot #(221, 10) dot22 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten22));
Dot #(230, 10) dot23 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten23));
Dot #(239, 10) dot24 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten24));
Dot #(13, 19) dot25 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten25));
Dot #(58, 19) dot26 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten26));
Dot #(112, 19) dot27 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten27));
Dot #(139, 19) dot28 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten28));
Dot #(194, 19) dot29 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten29));
Dot #(239, 19) dot30 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten30));
Dot #(58, 27) dot31 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten31));
Dot #(112, 27) dot32 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten32));
Dot #(139, 27) dot33 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten33));
Dot #(194, 27) dot34 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten34));
Dot #(13, 35) dot35 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten35));
Dot #(58, 35) dot36 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten36));
Dot #(112, 35) dot37 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten37));
Dot #(139, 35) dot38 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten38));
Dot #(194, 35) dot39 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten39));
Dot #(239, 35) dot40 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten40));
Dot #(13, 43) dot41 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten41));
Dot #(22, 43) dot42 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten42));
Dot #(31, 43) dot43 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten43));
Dot #(40, 43) dot44 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten44));
Dot #(49, 43) dot45 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten45));
Dot #(58, 43) dot46 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten46));
Dot #(67, 43) dot47 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten47));
Dot #(76, 43) dot48 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten48));
Dot #(85, 43) dot49 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten49));
Dot #(95, 43) dot50 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten50));
Dot #(104, 43) dot51 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten51));
Dot #(113, 43) dot52 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten52));
Dot #(122, 43) dot53 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten53));
Dot #(131, 43) dot54 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten54));
Dot #(140, 43) dot55 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten55));
Dot #(149, 43) dot56 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten56));
Dot #(158, 43) dot57 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten57));
Dot #(167, 43) dot58 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten58));
Dot #(176, 43) dot59 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten59));
Dot #(185, 43) dot60 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten60));
Dot #(194, 43) dot61 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten61));
Dot #(203, 43) dot62 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten62));
Dot #(212, 43) dot63 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten63));
Dot #(221, 43) dot64 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten64));
Dot #(230, 43) dot65 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten65));
Dot #(240, 43) dot66 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten66));
Dot #(13, 52) dot67 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten67));
Dot #(58, 52) dot68 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten68));
Dot #(85, 52) dot69 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten69));
Dot #(167, 52) dot70 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten70));
Dot #(194, 52) dot71 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten71));
Dot #(239, 52) dot72 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten72));
Dot #(13, 60) dot73 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten73));
Dot #(58, 60) dot74 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten74));
Dot #(85, 60) dot75 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten75));
Dot #(167, 60) dot76 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten76));
Dot #(194, 60) dot77 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten77));
Dot #(239, 60) dot78 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten78));
Dot #(13, 68) dot79 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten79));
Dot #(22, 68) dot80 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten80));
Dot #(31, 68) dot81 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten81));
Dot #(40, 68) dot82 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten82));
Dot #(49, 68) dot83 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten83));
Dot #(58, 68) dot84 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten84));
Dot #(85, 68) dot85 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten85));
Dot #(94, 68) dot86 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten86));
Dot #(103, 68) dot87 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten87));
Dot #(112, 68) dot88 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten88));
Dot #(139, 68) dot89 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten89));
Dot #(149, 68) dot90 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten90));
Dot #(158, 68) dot91 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten91));
Dot #(167, 68) dot92 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten92));
Dot #(194, 68) dot93 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten93));
Dot #(203, 68) dot94 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten94));
Dot #(212, 68) dot95 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten95));
Dot #(221, 68) dot96 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten96));
Dot #(230, 68) dot97 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten97));
Dot #(239, 68) dot98 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten98));
Dot #(58, 76) dot99 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten99));
Dot #(194, 76) dot100 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten100));
Dot #(58, 85) dot101 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten101));
Dot #(194, 85) dot102 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten102));
Dot #(58, 93) dot103 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten103));
Dot #(194, 93) dot104 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten104));
Dot #(58, 101) dot105 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten105));
Dot #(194, 101) dot106 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten106));
Dot #(58, 110) dot107 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten107));
Dot #(194, 110) dot108 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten108));
Dot #(58, 118) dot109 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten109));
Dot #(194, 118) dot110 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten110));
Dot #(58, 126) dot111 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten111));
Dot #(194, 126) dot112 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten112));
Dot #(58, 134) dot113 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten113));
Dot #(194, 134) dot114 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten114));
Dot #(58, 143) dot115 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten115));
Dot #(194, 143) dot116 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten116));
Dot #(58, 151) dot117 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten117));
Dot #(194, 151) dot118 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten118));
Dot #(58, 159) dot119 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten119));
Dot #(194, 159) dot120 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten120));
Dot #(13, 167) dot121 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten121));
Dot #(22, 167) dot122 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten122));
Dot #(31, 167) dot123 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten123));
Dot #(40, 167) dot124 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten124));
Dot #(49, 167) dot125 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten125));
Dot #(58, 167) dot126 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten126));
Dot #(67, 167) dot127 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten127));
Dot #(76, 167) dot128 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten128));
Dot #(85, 167) dot129 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten129));
Dot #(94, 167) dot130 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten130));
Dot #(103, 167) dot131 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten131));
Dot #(112, 167) dot132 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten132));
Dot #(140, 167) dot133 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten133));
Dot #(149, 167) dot134 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten134));
Dot #(158, 167) dot135 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten135));
Dot #(167, 167) dot136 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten136));
Dot #(176, 167) dot137 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten137));
Dot #(185, 167) dot138 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten138));
Dot #(194, 167) dot139 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten139));
Dot #(203, 167) dot140 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten140));
Dot #(212, 167) dot141 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten141));
Dot #(221, 167) dot142 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten142));
Dot #(230, 167) dot143 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten143));
Dot #(239, 167) dot144 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten144));
Dot #(13, 176) dot145 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten145));
Dot #(58, 176) dot146 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten146));
Dot #(112, 176) dot147 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten147));
Dot #(139, 176) dot148 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten148));
Dot #(194, 176) dot149 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten149));
Dot #(239, 176) dot150 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten150));
Dot #(13, 184) dot151 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten151));
Dot #(58, 184) dot152 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten152));
Dot #(112, 184) dot153 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten153));
Dot #(139, 184) dot154 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten154));
Dot #(194, 184) dot155 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten155));
Dot #(239, 184) dot156 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten156));
Dot #(22, 192) dot157 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten157));
Dot #(31, 192) dot158 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten158));
Dot #(58, 192) dot159 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten159));
Dot #(67, 192) dot160 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten160));
Dot #(76, 192) dot161 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten161));
Dot #(85, 192) dot162 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten162));
Dot #(94, 192) dot163 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten163));
Dot #(103, 192) dot164 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten164));
Dot #(112, 192) dot165 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten165));
Dot #(139, 192) dot166 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten166));
Dot #(148, 192) dot167 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten167));
Dot #(158, 192) dot168 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten168));
Dot #(167, 192) dot169 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten169));
Dot #(176, 192) dot170 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten170));
Dot #(185, 192) dot171 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten171));
Dot #(194, 192) dot172 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten172));
Dot #(221, 192) dot173 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten173));
Dot #(230, 192) dot174 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten174));
Dot #(31, 200) dot175 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten175));
Dot #(58, 200) dot176 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten176));
Dot #(85, 200) dot177 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten177));
Dot #(167, 200) dot178 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten178));
Dot #(194, 200) dot179 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten179));
Dot #(221, 200) dot180 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten180));
Dot #(31, 209) dot181 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten181));
Dot #(58, 209) dot182 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten182));
Dot #(85, 209) dot183 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten183));
Dot #(167, 209) dot184 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten184));
Dot #(194, 209) dot185 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten185));
Dot #(221, 209) dot186 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten186));
Dot #(13, 217) dot187 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten187));
Dot #(22, 217) dot188 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten188));
Dot #(31, 217) dot189 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten189));
Dot #(40, 217) dot190 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten190));
Dot #(49, 217) dot191 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten191));
Dot #(58, 217) dot192 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten192));
Dot #(85, 217) dot193 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten193));
Dot #(94, 217) dot194 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten194));
Dot #(103, 217) dot195 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten195));
Dot #(112, 217) dot196 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten196));
Dot #(139, 217) dot197 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten197));
Dot #(148, 217) dot198 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten198));
Dot #(158, 217) dot199 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten199));
Dot #(167, 217) dot200 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten200));
Dot #(194, 217) dot201 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten201));
Dot #(203, 217) dot202 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten202));
Dot #(212, 217) dot203 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten203));
Dot #(221, 217) dot204 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten204));
Dot #(230, 217) dot205 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten205));
Dot #(239, 217) dot206 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten206));
Dot #(13, 225) dot207 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten207));
Dot #(112, 225) dot208 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten208));
Dot #(139, 225) dot209 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten209));
Dot #(239, 225) dot210 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten210));
Dot #(13, 233) dot211 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten211));
Dot #(112, 233) dot212 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten212));
Dot #(140, 233) dot213 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten213));
Dot #(239, 233) dot214 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten214));
Dot #(13, 242) dot215 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten215));
Dot #(22, 242) dot216 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten216));
Dot #(31, 242) dot217 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten217));
Dot #(40, 242) dot218 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten218));
Dot #(49, 242) dot219 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten219));
Dot #(58, 242) dot220 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten220));
Dot #(67, 242) dot221 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten221));
Dot #(76, 242) dot222 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten222));
Dot #(85, 242) dot223 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten223));
Dot #(94, 242) dot224 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten224));
Dot #(103, 242) dot225 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten225));
Dot #(112, 242) dot226 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten226));
Dot #(121, 242) dot227 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten227));
Dot #(130, 242) dot228 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten228));
Dot #(139, 242) dot229 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten229));
Dot #(148, 242) dot230 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten230));
Dot #(158, 242) dot231 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten231));
Dot #(167, 242) dot232 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten232));
Dot #(176, 242) dot233 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten233));
Dot #(185, 242) dot234 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten234));
Dot #(194, 242) dot235 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten235));
Dot #(203, 242) dot236 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten236));
Dot #(212, 242) dot237 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten237));
Dot #(221, 242) dot238 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten238));
Dot #(230, 242) dot239 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten239));
Dot #(239, 242) dot240 (.Clk(VGA_VS), .Reset(Reset_h),.DrawX(DrawX), .DrawY(DrawY), .pac_mem_start_X(pac_mem_start_X), .pac_mem_start_Y(pac_mem_start_Y), .isEaten(isEaten240));



endmodule
